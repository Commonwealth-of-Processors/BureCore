`default_nettype none
module bure_stage_ex #()();
endmodule
`default_nettype wire
